module sll(out, a, b);



endmodule
