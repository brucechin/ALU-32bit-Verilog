module add_32()