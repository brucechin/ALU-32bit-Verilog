module alu_32(input [31:0] a, b,
              input [3:0] op,
              input [31:0] y,
              output carryout,
              output overflow,
              output zero,
              output [31:0] result);




endmodule