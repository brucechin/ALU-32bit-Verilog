module sll(a, movement, out);

output[31:0] out;
input[31:0] a;
input[4:0] movement;

assign out = 0;




endmodule
